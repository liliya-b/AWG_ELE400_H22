----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/30/2022 10:51:45 AM
-- Design Name: 
-- Module Name: Generator - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Generator is
    Port ( clk : in STD_LOGIC;
           reset : in STD_LOGIC;
           wave_type : in STD_LOGIC;
           dataout : out STD_LOGIC_VECTOR (7 downto 0));
end Generator;

architecture Wave_generator of Generator is

    CONSTANT TAILLE_ROM : positive := 40;
    TYPE romtype IS ARRAY (0 TO TAILLE_ROM) OF std_logic_vector(7 downto 0);
    
    signal i : integer := 0;

---- SINC WAVE WITH 40 SAMPLES----  
CONSTANT SincRom : romtype :=(
    0 =>    "00000001",  --0 : 1
    1 =>    "11110011",  --1 : -13
    2 =>    "11101000",  --2 : -24
    3 =>    "11100101",  --3 : -27
    4 =>    "11101100",  --4 : -20
    5 =>    "00000000",  --5 : 0
    6 =>    "00011110",  --6 : 30
    7 =>    "01000000",  --7 : 64
    8 =>    "01100000",  --8 : 96
    9 =>    "01110111",  --9 : 119
    10 =>   "01111111",  --10: 127
    11 =>   "01110111",  --11: 119
    12 =>   "01100000",  --12: 96
    13 =>   "01000000",  --13: 64
    14 =>   "00011110",  --14: 30
    15 =>   "00000000",  --15: 0
    16 =>   "11101100",  --16: -20
    17 =>   "11100101",  --17: -27
    18 =>   "11101000",  --18: -24
    19 =>   "11110011",  --19: -13
    20 =>   "00000000",  --20: 0
    21 =>   "00000000",  --21: 0
    22 =>   "00000000",  --22: 0
    23 =>   "00000000",  --23: 0
    24 =>   "00000000",  --24: 0
    25 =>   "00000000",  --25: 0
    26 =>   "00000000",  --26: 0
    27 =>   "00000000",  --27: 0
    28 =>   "00000000",  --28: 0
    29 =>   "00000000",  --29: 0
    30 =>   "00000000",  --30: 0
    31 =>   "00000000",  --31: 0
    32 =>   "00000000",  --32: 0
    33 =>   "00000000",  --33: 0
    34 =>   "00000000",  --34: 0
    35 =>   "00000000",  --35: 0
    36 =>   "00000000",  --36: 0
    37 =>   "00000000",  --37: 0
    38 =>   "00000000",  --38: 0
    39 =>   "00000000",  --39: 0
    40 =>   "00000000");  --40: 0

---- GAUSSIAN WAVE WITH 30 SAMPLES----  
CONSTANT GaussRom : romtype :=(
    0 =>    "00000010",  --0 : 2
    1 =>    "00000101",  --1 : 5
    2 =>    "00001000",  --2 : 8
    3 =>    "00001110",  --3 : 14
    4 =>    "00010110",  --4 : 22
    5 =>    "00100001",  --5 : 33
    6 =>    "00101111",  --6 : 47
    7 =>    "01000000",  --7 : 64
    8 =>    "01010010",  --8 : 82
    9 =>    "01100011",  --9 : 99
    10 =>   "01110010",  --10: 114
    11 =>   "01111100",  --11: 124
    12 =>   "01111111",  --12: 127
    13 =>   "01111100",  --13: 124
    14 =>   "01110010",  --14: 114
    15 =>   "01100011",  --15: 99
    16 =>   "01010010",  --16: 82
    17 =>   "01000000",  --17: 64
    18 =>   "00101111",  --18: 47
    19 =>   "00100001",  --19: 33
    20 =>   "00010110",  --20: 22
    21 =>   "00001110",  --21: 14
    22 =>   "00001000",  --22: 8
    23 =>   "00000101",  --23: 5
    24 =>   "00000010",  --24: 2
    25 =>   "00000000",  --25: 0
    26 =>   "00000000",  --26: 0
    27 =>   "00000000",  --27: 0
    28 =>   "00000000",  --28: 0
    29 =>   "00000000",  --29: 0
    30 =>   "00000000",  --30: 0
    31 =>   "00000000",  --31: 0
    32 =>   "00000000",  --32: 0
    33 =>   "00000000",  --33: 0
    34 =>   "00000000",  --34: 0
    35 =>   "00000000",  --35: 0
    36 =>   "00000000",  --36: 0
    37 =>   "00000000",  --37: 0
    38 =>   "00000000",  --38: 0
    39 =>   "00000000",  --39: 0
    40 =>   "00000000");  --40: 0

begin

PROCESS(clk)
    BEGIN
    
    IF(RISING_EDGE(clk)) THEN
    
        IF reset = '1' THEN
        
        i <= 0;
        
        ELSE
            
            IF wave_type = '1' then
            
             dataout <= GaussRom(i);
             
            ELSE 
            
             dataout <= SincRom(i);
        
            END IF;
            
            i<= i+1;
    
            IF(i = 40) THEN
            i<=0;
        
            END IF;
        END IF;
    END IF;
END PROCESS;

end Wave_generator;
