---- GAUSSIAN WAVE WITH 30 SAMPLES----  
CONSTANT GaussRom : romtype :=(
    0 =>    "01000000",  --0 : 64
    1 =>    "01001001",  --1 : 73
    2 =>    "01010010",  --2 : 82
    3 =>    "01011011",  --3 : 91
    4 =>    "01100011",  --4 : 99
    5 =>    "01101011",  --5 : 107
    6 =>    "01110010",  --6 : 114
    7 =>    "01110111",  --7 : 119
    8 =>    "01111100",  --8 : 124
    9 =>    "01111110",  --9 : 126
    10 =>   "01111111",  --10: 127
    11 =>   "01111110",  --11: 126
    12 =>   "01111100",  --12: 124
    13 =>   "01110111",  --13: 119
    14 =>   "01110010",  --14: 114
    15 =>   "01101011",  --15: 107
    16 =>   "01100011",  --16: 99
    17 =>   "01011011",  --17: 91
    18 =>   "01010010",  --18: 82
    19 =>   "01001001",  --19: 73
    20 =>   "01000000",  --20: 64
    21 =>   "00000000",  --21: 0
    22 =>   "00000000",  --22: 0
    23 =>   "00000000",  --23: 0
    24 =>   "00000000",  --24: 0
    25 =>   "00000000",  --25: 0
    26 =>   "00000000",  --26: 0
    27 =>   "00000000",  --27: 0
    28 =>   "00000000",  --28: 0
    29 =>   "00000000",  --29: 0
    30 =>   "00000000",  --30: 0
    31 =>   "00000000",  --31: 0
    32 =>   "00000000",  --32: 0
    33 =>   "00000000",  --33: 0
    34 =>   "00000000",  --34: 0
    35 =>   "00000000",  --35: 0
    36 =>   "00000000",  --36: 0
    37 =>   "00000000",  --37: 0
    38 =>   "00000000",  --38: 0
    39 =>   "00000000",  --39: 0
    40 =>   "00000000");  --40: 0